� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                             E~m~p~l~o~y~e~e~ ~N~a~m~e~ ~L~o~o~k~-~U~p~                                                                                                                                     Lpapsptp pNpapmpep                                                                   w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w                                         Fpiprpsptp pNpapmpep                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                