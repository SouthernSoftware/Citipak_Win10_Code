� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                   �������������������������������������������x                                     �O p p p p pE~m~p~l~o~y~e~e~ pQ~u~a~r~t~e~r~l~y~ ~W~a~g~e~ ~R~e~p~o~r~t~ p p p p p p�x                                     �O p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                     �O p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                     �O p p p pRpepppoprptp pupspipnpgp pQpupaprptpeprp:p           p p p p p p�                                     �O p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                     �O p p p p p p p p p p p p p p p p p p p pYpepaprp:p          p p p p p p p�                                     �O p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                     �O p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                     �O p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                     �O p p p p p p�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x p p p p p p�                                     �O p p p p p p��E~S~C~ ~Cpapnpcpeplp p���F~1~0~ ~Pprpopcpepspsp p� p p p p p p�                                     �O p p p p p p�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x p p p p p p�                                     ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  