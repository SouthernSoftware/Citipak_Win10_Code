� �  � �                      E{m{p{l{o{y{e{e{ {E{a{r{n{i{n{g{s{ {H{i{s{t{o{r{y{ {R{e{p{o{r{t{                      � REGION D CHILD CARE, INC.                                                       Employee Earnings History Report                                                Report D���������������������������������������������������������������x                 � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�         2       � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�          Trans D� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�   Hol      Reg E� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�oc Sec    RETIREM� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�ther 1   --------� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�---------10-31-19� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�  0.00      1,514� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p� 93.92         90� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p n p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�  0.00           � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�         10-31-19� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�  0.00      1,514� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p� 93.92         90� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�  0.00           � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�         10-28-19� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�  0.00      1,514� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p� 93.92         90� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�  0.00           ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�         09-27-1994        1784              Salaried       4.00       4.00       8.00      1,514.83       0.00       0.00       0.00       0.00   1,514.83      93.92    � ~F~1~ pHpeplppp p� pE~S~C~ pMpepnpup p� pF~5~ ~Pprpipnptp p� p p p p p p p p p� pH~o~m~e~ p� pE~n~d~ p� p~ p� p~ p� pP~g~U~p~ p� pP~g~D~n~ p� 