� �  �                                                                                                                                                                                                                                                                ������������������������������������������������x                                �                                              �                                �                                              �                                �                                              �                                �                                              �                                �                                              �                                �                                              �                                �                                              �                                ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�                                                                                                                                                                                                                                                                                                                                                                ������������������������������������������������x                                � �x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x �                                � ��F~1~ xHpeplppp�p��F~5~ xLpopopkpUppp�p��F~7~ pTpypppep�p��E~S~C~ xMpepnpup�p� �                                � �x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x �                                ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�                                                                                                                                                                                                                                                                                                                                                