� �  � � pFpepdpeprpaplp pTpapxp pTpapbplpep:p p pSpipnpgplpep p p p p p p p p p p p p p p p t t t t t t p p p p p p p p p p p p p p p pPpapgpep p1p popfp p2p p�                                                                                                  Employee Social Security %                                                      Employer Social Security %                                                      Social Security Max Wages $                                                     Employee Medicare %                                                             Employer Medicare %                                                             Medicare Max Wages $                                                            Std. Ded. Allow. Amount $                                                                                                                                                     T a x  T a b l e                                                  $ Amount           % Amount   On $ Amount Over                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        � ~F~1~ ~Hpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� pP~apgpepD~opwpnp p� p pPsasgsesUsps p p� 