� �  �                                                                                                                                                                                                                                                                                                                                                                                                                              ��������������������������������������������������x                               � p p p p p p p p p p pC~h~e~c~k~ ~P~r~i~n~t~i~n~g~ ~I~n~f~o~r~m~a~t~i~o~n~ p p p p p p p p p p p�x                               � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�x                               � p p p p p pSptpaprptpipnpgp pCphpepcpkp pNpupmpbpeprp:p                   p p�x                               � p p p p p p p p p p p p p p p p p p p p p p p p p p p p                   p p�x                               � p p p p p p p p p p p p pDpaptpep popfp pCphpepcpkpsp:p                   p p�x                               � p p p p p p p p p p p p p p p p p p p p p p p p p p p p                   p p�x                               � p p p p p p p p p p p p p p pPprpipnptpeprp pPpoprptp:p                   p p�x                               � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�x                               � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�x                               ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   � ~F~1~ ~Hpeplppp p p� p p p p p p p p p p p p p� pF~5~ ~ pAplpipgpnpmpepnptp pTpepsptp p� pF~1~0~ pPprpipnptp pCphpepcpkpsp p� pE~S~C~ ~Cpapnpcpeplp�p 