� �  ��� Ppapyprpoplplp pCpaplpcpuplpaptpipopnp p�p p p pEpmppplpopypepep:p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�p����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� p Earnings                                                                 p����� pRpepgp pEpaprpnpipnpgpsp p p p pOpTp pEpaprpnpipnpgpsp p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p����� p                                                                          p����� p Deductions                                                               p����� p p p pSpopcp pSpepcp p p p pMpepdpipcpaprpep p p p p pFpepdp pWp/pHp p p pSptpaptpep pWp/pHp p p p p p pRpeptpiprpep p p p p p p p p p p p p p p p p����� p                                                                          p����� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p����� p                                                                          p����� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p����� p                                                                          p����� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p��������������������������������������������������������������������������������������������������������������������������������������������������������������������� p   Gross Pay           Total Ded             Adv EIC           Net Pay    p����� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ~F~1~ ~Hpeplppp p p� pF~2~ pUpnpdpop p p p� pF~3~ ~Dpeplpeptpep p p� p p p p p ~ ~ ~ ~ ~ ~ ~ ~� pF~1~0~ pCpopnptpipnpupep p� pE~S~C~ ~Cpapnpcpeplp�p�