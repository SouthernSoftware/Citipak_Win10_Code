� �  � � pEpmppplpopypepep:p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�p                                                                                       1 Wages, tips other comp                2 Federal Income tax w/h                                                                                                3 Social Security wages                 4 Security Security w/h                                                                                                 5 Medicare wages and tips               6 Medicare tax w/h                                                                                                      7 Social Security tips                  8 Allocated tips                                                                                                        9 Advance EIC payment                  10 Dependent care benefits                                                                                              11 Nonqualified plans                   12 Benefits included in box 1                                                                                           13 See instrs. for box 13               14 Other                                                                                                                                                                                                15 Stat    Deceased  Pension   Legal      942    Subtotal  Deferred                 emp               plan      rep       emp                Comp                   [ ]      [ ]      [ ]       [ ]       [ ]      [ ]       [ ]                16 State  17 State wages, tips, etc     18 State Income taxes                                                                                                   19 Locality name    20 Local Wages      21 Local Income tax                                                                                                 � pF~1~ pHpeplppp p�p� p p p p p p p p�p� p p p p p p p p p�p� pE~s~c~ pMpepnpup p�p� p p p p p p p p p�p� p p p p p p p p p�p� pF~1~0~ pSpapvpep p�p 