� �  � � pSptpaptpep pTpapxp pTpapbplpep:p p pSpipnpgplpep p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p pPpapgpep p1p popfp p3p p�                                                                                                     Calc. Type (D or P)               ( )                                           Gross Wage Cut-Off Amt                                                          Min. Std. Adjust. Amt.                                                          Max. Std. Adjust. Amt.                                                          SUI %                                                                           SUI Max Wages                                                                   Std. Ded. Allow. Amount                                                                                                                                                      T a x   T a b l e                                                  $ Amount   % Amount      On $ Amount Over                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          � ~F~1~ ~Hpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� pP~apgpepD~opwpnp p� p pPsasgsesUsps p p� 