� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��������������������������������x                                                � pNpOp prpepcpoprpdpsp pipnp pEpmppplpopypepep pfpiplpep.p p�x                                                � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�x                                                � x x x x x x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x x x x x x x�x                                                � x x x x x x��������O~K~�p������� x x x x x x�x                                                � x x x x x x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x x x x x x x�x                                                ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       