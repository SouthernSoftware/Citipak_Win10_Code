� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ��������������������������������������������������x                              � p p p p p p p p p p pC~h~e~c~k~ ~P~r~i~n~t~i~n~g~ ~I~n~f~o~r~m~a~t~i~o~n~ p p p p p p p p p p p�x                              �  p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p �x                              �        Sptpaprptpipnpgp pCphpepcpkp pNpupmpbpeprp p:p             p p p p �x                              �  p p p p p p p p p p p p p pDpaptpep popfp pCphpepcpkpsp p:p             p p p p �x                              �  p p p p p p p p p p p p p p p pPprpipnptpeprp pPpoprptp p:p               p p �x                              �  p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p �x                              �   �x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x x p �x                              �  p p�x� ~F~1~ pHpeplppp p p p� pE~S~C~ pCpapnpcpeplp p� pF~1~0~ pCpopnptpipnpupep�p�x x p �x                              �  p p�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x p p �x                              ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 