� �  �                                                                                                                                                                This procedure removes the cleared checks from the outstanding                  check file.                                                                                                                                                     Press any key to continue or Esc to cancel.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     