� �  �                                                                                   p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p      p p p p p p p p p p p p p p p p p p p p p p pE~m~p~l~o~y~e~e~ ~Y~e~a~r~ ~t~o~ ~D~a~t~e~ ~T~o~t~a~l~s~ ~ p p p p p p p p p p p p p p p p p p p p p p p      p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p      p Gross - Net - EIC - Other Earnings                                       p      pRpepgp pEpaprpnpipnpgpsp p p p pOpTp pEpaprpnpipnpgpsp p p p p p p p p pEpaprpnp p1p p p p p p p p p pEpaprpnp p2p p p p p p p p p pEpaprpnp p3p p p      p p p p p9p,p1p0p0p.p0p0p p p p p p p p7p,p9p9p0p.p0p0p p p p p p p p6p,p9p9p0p.p0p0p p p p p p p p5p,p9p9p0p.p0p0p p p p p p p p4p,p9p9p0p.p0p0p p p       p p p p p pNpeptp pPpapyp p p p p p p p pApdpvp pEpIpCp p p p p pTpoptpaplp pEpaprpnp p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p      p p p p p6p,p9p9p0p.p0p0p p p p p p p p5p,p9p9p0p.p0p0p p p p p p p p4p,p9p9p0p.p0p0p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p      p p p pGprpopspsp pPpapyp p p p p p pFpepdp pGprpopspsp p p p pSptpaptpep pGprpopspsp p p p p p pMpepdp pGprpopspsp p p p p p pSpopcp pGprpopspsp p p      p p p p p1p,p0p0p0p.p0p0p p p p p p p p1p,p0p0p0p.p0p0p p p p p p p p1p,p0p0p0p.p0p0p p p p p p p p1p,p0p0p0p.p0p0p p p p p p p p1p,p0p0p0p.p0p0p p p      p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p      p Deductions - Taxes - Retirement                                          p      p p p p pSpopcp pSpepcp p p p pMpepdpipcpaprpep p p p p pFpepdp pWp/pHp p p pSptpaptpep pWp/pHp p p p p p pRpeptpiprpep p p pTpoptpaplp pDpepdp p p p      p p p9p9p,p9p9p9p.p0p2p p p p9p9p,p9p9p9p.p9p9p p p p9p9p,p6p2p0p.p1p7p p p p9p9p,p8p2p0p.p0p7p p p p9p9p,p7p4p8p.p6p0p p p p9p9p,p9p9p0p.p0p0p p p p      p p p pCpapfpep pIpnpsp p p pIpnpspuprpapnpcpep p p p p p p pOptphpeprp p p p p p p pOptphpeprp p p p p p p pOptphpeprp p p p p p p pOptphpeprp p p p      p p p p9p,p1p0p0p.p0p0p p p p p8p,p9p9p0p.p0p0p p p p p7p,p9p9p0p.p0p0p p p p p6p,p9p9p0p.p0p0p p p p p5p,p9p9p0p.p0p0p p p p p4p,p9p9p0p.p0p0p p p p      p p p p p p pOptphpeprp p p p p p p p p pYpopup p p p p p p p p pCpapnp p p p p p pCphpapnpgpep p p p p p p pTphpepspep p p p p p p pOptphpeprp p p p      p p p p9p,p1p0p0p.p0p0p p p p p8p,p9p9p0p.p0p0p p p p p7p,p9p9p0p.p0p0p p p p p6p,p9p9p0p.p0p0p p p p p5p,p9p9p0p.p0p0p p p p p4p,p9p9p0p.p0p0p p p p      p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p      p p p p p p p p p p p p p p p p p p�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q p p p p p p p p p p p p p p p p p p p p p      p p p p p p p p p p p p p p p p p p �q        � pO~K~ ~ pCpopnptpipnpupep p�           p p p p p p p p p p p p p p p p p p p p p      p p p p p p p p p p p p p p p p p p�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q�q p p p p p p p p p p p p p p p p p p p p p                                                                                                                                                                   