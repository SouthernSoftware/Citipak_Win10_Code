� �  � � pEpmppplpopypepep pLpepapvpep pBpepnpepfpiptp pMpapipnptpepnpapnpcpep p p p p p p p p p p p p p p p p p p p p p p p p p p p p pPpapgpep p1p popfp p1p p�                                                                                        Employee Leave File Options                                                                                                                                         Vacation Benefit             Maximum Accrued                                             Years of Service                                                                Over-       But not over-      Hours Earned                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       Sick Leave                  Maximum Accrued                                             Years of Service                                                                Over-       But not over-      Hours Earned                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            � pF~1~ pHpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� p p p p p p p p p p p� p p p p p p p p p� 