� �  �                                                                                                                                                                                                                                                                �������������������������������������������������x                               �  p p p p p pE~m~p~l~o~y~e~e~ ~E~a~r~n~i~n~g~s~ ~H~i~s~t~o~r~y~ ~R~e~p~o~r~t~ p p p p p p p p�x                               �  p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p �x                               �  p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p �x                               �  p p p p p pFpiprpsptp pEpmppplpopypepep pNpop:p                      �x                               �  p p p p p p p p p p p p p p p p p p p p p p p p                      �x                               �  p p p p p p pLpapsptp pEpmppplpopypepep pNpop:p                      �x                               �  p p p p p p p p p p p p p p p p p p p p p p p p                      �x                               �  p p p p p p p p p p p p pSptpaprptp pDpaptpep:p                      �x                               �  p p p p p p p p p p p p p p p p p p p p p p p p                      �x                               �  p p p p p p p p p p p pEpnpdpipnpgp pDpaptpep:p                      �x                               �                                       p p p p p p p p �x                               �         �x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x       x p �x                               �         ��E~S~C~ ~Cpapnpcpeplp p���F~1~0~ ~Pprpopcpepspsp p�       x p �x                               �         �x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x       p p �x                               ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               