� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�O�x                                         � N N N NINnNvNaNlNiNdN NSNtNaNrNtNiNnNgN NCNhNeNcNkN NNNuNmNbNeNrN N N N N�                                         � N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N�                                         � N N NPKlKeKaKsKeK KEKnKtKeKrK KaK KNKEKWK NCKhKeKcKkK KNKuKmKbKeKrK K N N�                                         � N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N N�                                         � N N N N N N N N N N N N N�H�H�H�H�H�H�H�H�H�H N N N N N N N N N N N N N N�                                         � N N N N N N N N N N N N N�� ~ ~O~K~ ~ ~�p� N N N N N N N N N N N N N N�                                         � N N N N N N N N N N N N N�H�H�H�H�H�H�H�H�H�H N N N N N N N N N N N N N N�                                         ��H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�H�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     