� �  � � pMpapnpupaplp pTprpapnpspapcptpipopnp pEpnptprpyp p:p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                                                                   Period Beg:           End:               Voluntary Deductions                   Check Date:            No:               Description             Amount         Hours Worked:                                                                   Sick Hours:                                                                     Vacation Hours:                                                                 Comp Hrs:                                                                       Holiday Hrs:                                                                    OT Hrs Paid:                                                                    Wage Distributions                                                              G/L Acct Number        Amount                                                   1)                                                                              2)                                                                              3)                                                                              4)                                                                              Gross Pay:                               Total Vol Deductions:                  REG:             OT:                     Earned Income Credit:                      Federal Tax W/H:                           Net Pay:                               State Tax W/H:                     Federal Gross:                         Social Security W/H:                       State Gross:                                Medicare W/H:                      Social Gross:                              Retirement W/H:                    Medicare Gross:                                                                      c                                 � ~F~1~ ~Hpeplppp p p� p p p p p p p p p p p� pF~3~ ~Dpeplpeptpep p p� p p p p p ~ ~ ~ ~ ~ ~ ~ ~� pF~1~0~ pCpopnptpipnpupep p� pE~S~C~ ~Cpapnpcpeplp�p 