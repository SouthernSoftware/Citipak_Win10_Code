� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                            E~m~p~l~o~y~e~e~ ~N~u~m~b~e~r~ ~L~o~o~k~-~U~p~                                                                                                                                w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w                                        Epmppplpopypepep pNpop                                                                   w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   