� �  � � pEpmppplpopypeprp pIpnpfpoprpmpaptpipopnp pFpiplpep p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                                                                                                                                                                                                                                                                                                                                    Employer Name                                                                       Attention                                                                         Address                                                                         Address                                                                            City                                                                           State                                                                             Zip                                                                      Fed Tax ID                                                                    State Tax ID                                                                    Ret Sys ID-G                                                                    Ret Sys ID-L                                                                                                                                                 ESC Report Type                                                               Taxable Wage Base                                                                                                                                                    BB&T Center#                                                                          Batch#                                                                                                                                                                                                                 � ~F~1~ ~Hpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� p p p p p p p p p p� p p p p p p p p p p� 