� �  � � pEpmppplpopypepep pMpapipnptpepnpapnpcpep:p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p pPpapgpep p1p popfp p3p p�                                                                                   Employee Information                                                                                                                                                 Number                          Soc Sec No                                   Last Name                          First Name                                     Address                                                                         Address                                                                            City                               State          Zip                      Birthdate                              Gender         Race                     Ret Number                            Ret Type                                  DD Acct No                                                                                                                                                                                                                                     Job Description                                                                                                                                                       Title                                         W/C Code                         Status             Benefit Pct                 Pay Type                      Frequency                    Rate                O/T  Rate                      Hire Date             Next Review                Term Date                                                                                                                                                                                                                                                                                                                                                   � ~F~1~ ~Hpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� pF~7~ pYp-pTp-pDp p� pP~apgpepD~opwpnp p� p pPsasgsesUsps p p� 