� �  � � pSpypsptpepmp pCpopnptprpoplp pFpiplpep p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                                                                                                                                                        Imprest Payroll Acct                                                               Imprest Cash Acct                                                          Imprest Wages Pay Acct                                                          Print PR Deposit Check                                                             Imprest Vendor Code                                                                                                                                             Federal W/H Acct No                                                               State W/H Acct No                                                             Soc Sec W/H Acct No                                                            Medicare W/H Acct No                                                          Retirement W/H Acct No                                                                                                                                         Calculate Expense Match                                                                Soc Sec Exp Code                                                               Medicare Exp Code                                                             Retirement Exp Code                                                             Due to Account Code                                                           Due From Account Code                                                                Interface to G/L                                                                                                                                                                                                                      � ~F~1~ ~Hpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� p p p p p p p p p p� p p p p p p p p p p� 