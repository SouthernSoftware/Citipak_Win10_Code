� �  ��� Ppapyprpoplplp pTprpapnpspapcptpipopnpsp�p pEpmppplpopypepep:p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�p������������������������������������������������������������������������������������� p Hours this Period                    Distribution                     p�������� p p p p p p pRpepgpuplpaprp pHpopuprpsp pWpoprpkpepdp          p p ?G?/?L? ?A?c?c?o?u?n?t?#? ? ?�? ?R?e?g? ?H?r?s?�? ?O?/?T? ?H?r?s? p�������� p p p p p p p pVpapcpaptpipopnp pHpopuprpsp pUpspepdp          p py              �        �         p�������� p p p p p p p p p p p pSpipcpkp pHpopuprpsp pUpspepdp          p py              �        �         p�������� p p p p p p p p pHpoplpipdpapyp pHpopuprpsp pUpspepdp          p py              �        �         p�������� p p p p p p p p p p p pCpopmppp pHpopuprpsp pPpapipdp          p py              �        �         p�������� p p pTpoptpaplp pRpepgpuplpaprp pHpopuprpsp pPpapipdp ~ ~ ~ ~ ~ ~ ~ ~ ~ p py              �        �         p�������� p p p p p pOpvpeprptpipmpep pHpopuprpsp pWpoprpkpepdp          p py              �        �         p�������� p p p p p p p pOpvpeprptpipmpep pHpopuprpsp pPpapipdp ~ ~ ~ ~ ~ ~ ~ ~ ~ p py              �        �         p�������� p p p p pOpvpeprptpipmpep pHpopuprpsp ptpop pCpopmppp          p py              �        �         p�������� p p p p p p p p p p p p p p p p p p p p p p p p p p p          p pyTpoptpaplpsp p p p p p p p p� ~ ~ ~ ~ ~ ~ ~ ~� ~ ~ ~ ~ ~ ~ ~ ~ p�������� p Additional Earnings                  Addit'l Earnings Distribution    p�������� p p p p p p p p p p p p p p p p p p p p p p p p p p.p          p p ?G?/?L? ?A?c?c?o?u?n?t?#? ? ? ? ? ? ?�? ? ? ? ? ? ? ?A?m?o?u?n?t? p�������� p p p p p p p p p p p p p p p p p p p p p p p p p p.p          p py                  �              p�������� p p p p p p p p p p p p p p p p p p p p p p p p p p.p          p py                  �              p�������� p p p p p p p p p p p p p p p p p p p p p p p p p p p          p py                  �              p�������� p p p p p p p p p p p p p p p p p p p p p p p p p p p          p py                  �              p�������� p p p p p p p p p p p p p p p p p p p p p p p p p p p          p py                  �              p�������� p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p py                  �              p�������� pTpoptpaplp pApdpdp'plp pEpaprpnpipnpgpsp p.p.p.p.p.p ~ ~ ~ ~ ~ ~ ~ ~ ~ p pyTpoptpaplpsp p p p p p p p p p p p p� ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ ~ p���������������������������������������������������������������������������������������������������������������������������������������������������������������������� ~F~1~ ~Hpeplppp p p� pF~2~ pUpnpdpop p p p� pF~3~ ~Dpeplpeptpep p p� p p p p p ~ ~ ~ ~ ~ ~ ~ ~� pF~1~0~ pCpopnptpipnpupep p� pE~S~C~ ~Cpapnpcpeplp�p�