� �  ��� Epdpiptp p/p pVpipepwp pEpmppplpopypepep pIpnpfpoprpmpaptpipopnp p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�x������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ~F~1~ ~Hpeplppp p� pF~5~ pSpepaprpcphp p� p p p p p p p p p� pF~7~ pNpapmpep p p p� p p p p p p p p p p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p�x�