� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������������������������������������������������x                                � p p ~ ~ ~ ~ ~ ~ ~ ~ ~ pE~m~p~l~o~y~e~e~ ~N~a~m~e~ ~L~o~o~k~-~U~p~ p p p p p p p p p p p p p�                                � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                � p p pLpapsptp pNpapmpep                                  p�                                � p p p p p p p p p p p p                                  p�                                � p pFpiprpsptp pNpapmpep                                  p�                                � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                � p�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x p�                                � p���F~1~ xHpeplppp�p������F~5~ xLpopopkpUppp�p������E~S~C~ xMpepnpup�p�� p�                                � p�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x p�                                ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               