� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ������������������������������������x                                                � p pLpapsptp pApcpcprpupaplp pDpaptpep:p p1p2p/p1p3p/p1p9p9p4p w p p�x                                                � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p w p p�x                                                � p p p p pApcpcprpupep pTphprpopupgphp:p p p p p p p p p p p p w p p�x                                                � p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�x                                                � x x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x x x�x                                                � x x����E~S~C~ ~Cpapnpcpeplp�p��F~1~0~ ~Upppdpaptpep�p�� x x�x                                                � x x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x x x�x                                                ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           