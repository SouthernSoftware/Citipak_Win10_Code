� �  � � pWp-p2p pEpxptprpapcptpipopnp pSpeptpuppp p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�p                                                                                                                                                                                                                 Amount in                                Deduction        Check box               Box            Code                                                                                                    Retirement                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              � pF~1~ pHpeplppp p�p� p p p p p p p p�p� p p p p p p p p p�p� pE~s~c~ pMpepnpup p�p� p p p p p p p p p�p� p p p p p p p p p�p� pF~1~0~ pSpapvpep p�p 