� �  � � pEpmppplpopypepep pMpapipnptpepnpapnpcpep:p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p pPpapgpep p3p popfp p3p p�                                                                                   Default Earning Codes                                                              Description           Account Number     Earnings                                                                                                                                                                                                                                                                                                                                                         Wage Distribution                                                                              Account Number         Default Distribution                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Benefit Schedule              Earned           Used       Balance                            Vacation                                                                        Sick Leave                                                                      Comp Time                                                                                                                                         � ~F~1~ ~Hpeplppp p� pF~4~ pHpipsptpoprpyp p� pF~7~ pYp-pTp-pDp p� p pP~apgpepD~np p p� pP~apgpepU~pp p p� pF~1~0~ pSpapvpep p� pE~S~C~ ~Mpepnpup p� 