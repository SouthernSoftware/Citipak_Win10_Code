� �  � � pPprpipnptpeprp pSpeptpuppp p&p pCpopnpfpipgpuprpaptpipopnp p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p�                                                                                                                                                                                                                                                                                                                                                    Employee Data File                                                            Active Employee List                                                        Terminated Employee List                                                       Employee Earnings History                                                                Quarterly Report                                                        Payroll Deductions Taken                                                                      ESC Report                                                            Leave Benefit Report                                                          YTD Wage Distributions                                                              Retirement Reports                                                         Supplemental Retirement                                                                                                                                 Payroll Register & Distribution                                                             GL Interface Report                                                                  Payroll Checks                                                          Payroll Check Register                                                                                                                                                                                                                                                                                            � ~F~1~ ~Hpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� p p p p p p p p p p� p p p p p p p p p p� 