� �  � � pEpmppplpopypepep pMpapipnptpepnpapnpcpep:p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p pPpapgpep p2p popfp p3p p�                                                                                   Tax Withholding                                                                                         Fixed                                                              Exempt  Amt/Pct  Figure   Status   # Allowances   Addit W/H Amt       Federal                                                                         State                                                                           Social Security Exempt?         Medicare Exempt?       EIC Code                                                                                                Misc Deductions                                                                    Description             Amt/Pct       Withhold     Inc O/T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � ~F~1~ ~Hpeplppp p� pF~4~ pHpipsptpoprpyp p� pF~7~ pYp-pTp-pDp p� p pP~apgpepD~np p p� pP~apgpepU~pp p p� pF~1~0~ pSpapvpep p� pE~S~C~ ~Mpepnpup p� 