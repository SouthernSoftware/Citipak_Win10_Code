� �  � � pEpaprpnpipnpgpsp pCpopdpep pMpapipnptpepnpapnpcpep p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p pPpapgpep p1p popfp p1p p�                                                                                        Earnings File Options                                                                                                                                                                                                                                   Description             Withhold on Earnings                                                    FWT     SWT     SOC     MED    RET                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          � pF~1~ pHpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� pF~8~ pRpepmpopvpep p� p p p p p p p p p� 