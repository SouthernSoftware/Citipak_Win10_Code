� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ���������������������������������������������������x                             � p p p p p p p p p p p p p p p p p p p p p p p p p�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x p p�x                             � p pSptpaprptp:p p p p p p p p p p p p p p p p p p�x�F~5~ ~ pAplpipgpnpmpepnptp pTpepsptp�p�x p p�x                             � p p pDpaptpep:p p p p p p p p p p p p p p p p p p�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x p p�x                             � p p p p p p p p p p p p p p p p p p p p p p p p p�x�F~1~0~ pPprpipnptp pCphpepcpkpsp p p�p�x p p�x                             � p p p p p p p p p p p p p p p p p p p p p p p p p�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x p p�x                             � p p p pRpepapdpyp ptpop pPprpipnptp p p p p p p p�x�E~S~C~ pApbpoprptp p p p p p p p p p�p�x p p�x                             � p p p p p p pCphpepcpkpsp?p p p p p p p p p p p p�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x p p�x                             ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               