� �  � � pEpaprpnpepdp pIpnpcpopmpep pCprpepdpiptp pTpapbplpep:p pMpaprprpipepdp pwpiptphp pSpppopupspep pCpeprptpipfpipcpaptpep p p p p p p p p p p p p p p p p�                                                                                                                                                                                                                                                                                                                                         Annualized Wages                                                                (Before withholding                                                             allowances)                                                                                                     Amt of                Of wages in                 Over-       But not over-     Payment       Less      excess of                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        � ~F~1~ ~Hpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� pP~apgpepD~opwpnp p� p pPsasgsesUsps p p� 