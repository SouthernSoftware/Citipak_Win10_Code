� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                �O�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�_�x                                  �O _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _�                                  �O _ _ _ _ _ _ _ _P^a^y^r^o^l^l^ ^D^e^m^o^n^s^t^r^a^t^i^o^n^ ^V^e^r^s^i^o^n^ _ _ _ _ _ _ _�                                  �O _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _�                                  �O _ _ _Y_o_u_ _m_a_y_ _O_N_L_Y_ _e_d_i_t_ _a_n_ _e_x_i_s_t_i_n_g_ _E_m_p_l_o_y_e_e_._ _ _�                                  �O _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _�                                  �O _ _ _ _P_l_e_a_s_e_ _c_o_n_t_a_c_t_ _S_o_u_t_h_e_r_n_ _S_o_f_t_W_a_r_e_ _f_o_r_ _ _ _ _�                                  �O _ _ _ _a_d_d_i_t_i_o_n_a_l_ _i_n_f_o_r_m_a_t_i_o_n_._ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _�                                  �O _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _�                                  �O _ _ _ _ _ _ _ _ _ _ _ _ _ _1^-^8^0^0^-^8^4^2^-^8^1^9^0^ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _�                                  �O _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _�                                  �O _ _ _ _ _ _ _ _ _P^r^e^s^s^ ^a^n^y^ ^K^e^y^ ^t^o^ ^c^o^n^t^i^n^u^e^.^ _ _ _ _ _ _ _ _ _�                                  �O _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _ _�                                  ��X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�X�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  