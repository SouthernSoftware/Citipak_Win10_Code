� �  � � pRpeptpiprpepmpepnptp pFpiplpep pMpapipnptpepnpapnpcpep p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p pPpapgpep p1p popfp p1p p�                                                                                        Retirement File Options                                                                                                                                                                                                                                                      Withholding    Matching    Include                  Type Description            Rate           Rate        Overtime                                                                                                  1                                                                               2                                                                               3                                                                               4                                                                               5                                                                               6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       � pF~1~ pHpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� pF~8~ pRpepmpopvpep p� p p p p p p p p p� 