� �  �  P pPpapyprpoplp pTprpapnpspapcptpipopnpsp p�p pLpapsptp pEpmppplpopypep pEpnptpeprpepdp p:p p����@� ?T?r?a?n?s?a?c?t?i?o?n? ?E?n?t?r?y? ?/? ?E?d?i?t? ? �. p�� pEpmppp pNpupmpbpeprp! p��. p��. p��/�������-� pFp1p-pHpeplppp pEpSpCp-pApbpoprptp pFp1p0p-pCpopnptpipnpupep+ p������������������������������������������������������������������x��������� p p p p p p p p p p p p p p p p p p p p ~P~r~o~c~e~s~s~i~n~g~ ~D~a~t~e~s~ ~/~ ~O~p~t~i~o~n~s~ ~ p p p p p p p p p p p p p p p p p p p p p p�x���������                                                                      �x��������� Ppapyp pPpeprpipopdp pBpepgpipnpnpipnpgp pDpaptpep                Epnpdpipnpgp pDpaptpep                 �x���������                                                                      �x��������� S~e~t~ ~P~a~y~r~o~l~l~ ~w~i~t~h~ ~D~e~f~a~u~l~t~s~?~ (p )p p p p p p p p p p p p p p p p                        �x��������� Epmppplpopypepepsp ptpop pPpapyp:p p                                                   �x���������  p p p p p p p p p pWpepepkplpyp p p(p )p p p p p p p p p p p pMpopnptphplpyp p p(p )p            pApnpnpupaplpyp p p(p )p �x���������  p p p p p p pBpip-pWpepepkplpyp p p(p )p p p p p p p p p pQpupaprptpeprplpyp p p(p )p                         �x���������  p p p pSpepmpip-pMpopnptphplpyp p p(p )p p p p p p pSpepmpip-pApnpnpupaplpyp p p(p )p                         �x���������                       p p p p p p p p p p p p p p p p p p p p p p p p                        �x��������� D~e~d~u~c~t~i~o~n~s~ ~t~o~ ~t~a~k~e~ ~                                                  �x���������   1p)p p p p p p p p p p p p p p p(p )p p p p p5p)p p p p p p p p p p p p p p p(p )p p p p p p9p)p p p p p p p p p p p p p p p(p )p p�x���������   2p)p p p p p p p p p p p p p p p(p )p p p p p6p)p p p p p p p p p p p p p p p(p )p p p p p1p0p)p p p p p p p p p p p p p p p(p )p p�x���������   3p)p p p p p p p p p p p p p p p(p )p p p p p7p)p p p p p p p p p p p p p p p(p )p p p p p1p1p)p p p p p p p p p p p p p p p(p )p �x���������   4p)p p p p p p p p p p p p p p p(p )p p p p p8p)p p p p p p p p p p p p p p p(p )p p p p p1p2p)p p p p p p p p p p p p p p p(p )p �x���������                                                                      �x��������� A~d~d~i~t~i~o~n~a~l~ ~E~a~r~n~i~n~g~s~ ~A~c~c~o~u~n~t~s~ ~t~o~ ~u~s~e~                                  �x���������   1p)p p p p p p p p p p p p p p p(p )p p p p p2p)p p p p p p p p p p p p p p p(p )p p p p p p3p)p p p p p p p p p p p p p p p(p )p �x����������x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�������������������������������������������������������������������������������������������������������������������������������������������������������������������� pFp1p-pHpeplppp p p pEpSpCp-pApbpoprptp p p p pFp1p0p-pCpopnptpipnpupep p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p