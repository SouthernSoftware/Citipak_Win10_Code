� �  � � pDpepdpupcptpipopnp pCpopdpep pMpapipnptpepnpapnpcpep p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p p pPpapgpep p1p popfp p1p p�                                                                                        Deduction File Options                                                                                                                                                                                Withholding Exemptions                       #  Description   Liab Acct #     FWT     SWT     SOC     MED                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            � pF~1~ pHpeplppp p p� pF~1~0~ pSpapvpep p� p p p p p p p p p p� pE~S~C~ ~Mpepnpup p� p p p p p p p p p p� pF~8~ pRpepmpopvpep p� p p p p p p p p p� 