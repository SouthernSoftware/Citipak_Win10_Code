� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ����������������������������x                                                    � p p p p p p p pSpcpapnpnpipnpgp.p.p.p p p p p p p p�x                                                    � x p p p p p p p p p p p x x x x x x x x x x x x x x�x                                                    � x x p p p p p p p p pcpopmppplpeptpepdp.p p x x x x�x                                                    ��x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x�x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         